package riscv_pkg;
	import uvm_pkg::*;

	`include "riscv_sequencer.sv"
	`include "riscv_monitor.sv"
	`include "riscv_driver.sv"
	`include "riscv_agent.sv"
	`include "riscv_scoreboard.sv"
	`include "riscv_config.sv"
	`include "riscv_env.sv"
	`include "riscv_test.sv"
endpackage: riscv_pkg
