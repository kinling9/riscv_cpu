module riscv_hazard(

);
// 该模块对于冒险信号进行检测，并生成对应的调度信号
endmodule