interface control_if;
  logic clk;
  logic rst_n;
  logic [31:0] i_boot_addr;
endinterface: control_if