class riscv_configuration extends uvm_object;
	`uvm_object_utils(riscv_configuration)

	function new(string name = "");
		super.new(name);
	endfunction: new
endclass: riscv_configuration
